module logic(

    );
endmodule
