module ADD(
    input 

    );
endmodule

module SUB(
    input wire

    );
endmodule

module SHL(
    input wire

    );
endmodule

module SHR(
    input wire

    );
endmodule

module CMP(
    input wire

    );
endmodule

module AND(
    input wire

    );
endmodule

module OR(
    input wire

    );
endmodule

module XOR(
    input wire

    );
endmodule

module NAND(
    input wire

    );
endmodule

module NOR(
    input wire

    );
endmodule

module XNOR(
    input wire

    );
endmodule

module INV(
    input wire

    );
endmodule

module NEG(
    input wire

    );
endmodule

module STO(
    input wire

    );
endmodule

module SWP(
    input wire

    );
endmodule

module LOAD(
    input wire

    );
endmodule




